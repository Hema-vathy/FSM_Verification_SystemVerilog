//////////////*************INTERFACE FILE - CONTAIN ALL THE SIGNAL NEEDED FOR THE VERIFICATION*************//////////////
interface signal;
  logic clock;
  logic reset;
  logic sequence_in;
  logic detector_out;
  logic sequence_q[$];
endinterface
