/////////////*************PACKAGE CONTAINING FILES*************/////////////
package pkg;
`include "clk_gen.sv"
`include "stimuli.sv"
`include "rst_gen.sv"
`include "reset_test.sv"
`include "comparison_test.sv"
`include "run_test.sv"
endpackage
